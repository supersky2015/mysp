test array
vin1 1 0 10.0 ac 1.0 sin(0 1 10 )
vin2 2 0 10.0 ac 1.0 sin(0 1 10 -0.03333333333)
vin3 3 0 10.0 ac 1.0 sin(0 1 10 -0.06666666666)
R1 1 0 2
r2 2 0 2
r3 3 0 2
.tran 100u 0.2 uic